LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux8_32bits IS
PORT(
	DIn0 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	DIn1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	DIn2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	DIn3 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	DIn4 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	DIn5 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	DIn6 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	DIn7 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	ctrl : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	Dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
);
END mux8_32bits;

ARCHITECTURE mux8_32bits_behavior OF mux8_32bits IS
BEGIN

WITH ctrl SELECT Dout <= DIn0 WHEN "000",
		DIn1 WHEN "001",
		DIn2 WHEN "010",
		DIn3 WHEN "011",
		DIn4 WHEN "100",
		DIn5 WHEN "101",
		DIn6 WHEN "110",
		DIn7 WHEN OTHERS;

END mux8_32bits_behavior;
