LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux8_32bits IS
PORT(
	Din0 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	Din1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	Din2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	Din3 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	Din4 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	Din5 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	Din6 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	Din7 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
	ctrl : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
	Dout : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
);
END mux8_32bits;

ARCHITECTURE mux8_32bits_behavior OF mux8_32bits IS
BEGIN

WITH ctrl SELECT Dout <= DIn0 WHEN "000",
		Din1 WHEN "001",
		Din2 WHEN "010",
		Din3 WHEN "011",
		Din4 WHEN "100",
		Din5 WHEN "101",
		Din6 WHEN "110",
		Din7 WHEN OTHERS;

END mux8_32bits_behavior;